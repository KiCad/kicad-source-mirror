.title KiCad schematic
.include "chirp.lib.spice"
.save all
.probe alli
.tran 10u 100m

R1 /out Net-_V1-E2_ 10k 
XV1 /out Net-_V1-E2_ chirp bf=1k ef=3k bt=30m et=70m 
.end
