.title KiCad schematic
.include "opamp.lib"
.save all
.probe alli
.tran 10u 10m

R1 GND Net-_U1--_ 10k 
R2 Net-_U1--_ /out 10k 
V3 GND Net-_U1-V-_ ( 5 ) 
VSIN1 /in GND SIN( 0 100m 1k ) 
V2 Net-_U1-V+_ GND ( 5 ) 
XU1 /in Net-_U1--_ Net-_U1-V+_ Net-_U1-V-_ /out uopamp_lvl2 
.end
