*
* fets.lib.spice
*

* All parameter values are made up and physically nonsensical.

.model _0_NJF_SHICHMANHODGES njf (level=1
+ VTO=000.000E+07
+ BETA=100.001E+07
+ LAMBDA=200.002E+07
+ RD=300.003E+07
+ RS=400.004E+07
+ CGS=500.005E+07
+ CGD=600.006E+07
+ PB=700.007E+07
+ IS=800.008E+07
+ FC=900.009E+07
+)

.model _1_PJF_SHICHMANHODGES pjf (level=1
+ VTO=000.000E+07
+ BETA=100.001E+07
+ LAMBDA=200.002E+07
+ RD=300.003E+07
+ RS=400.004E+07
+ CGS=500.005E+07
+ CGD=600.006E+07
+ PB=700.007E+07
+ IS=800.008E+07
+ FC=900.009E+07
+)

.model _2_NJF_PARKERSKELLERN njf (level=2
+ VBI=000.000E+07;;;
+ AF=100.001E+07
+ BETA=200.002E+07
+ CDS=300.003E+07
+ CGD=400.004E+07
+ CGS=500.005E+07
+ DELTA=600.006E+07
+ HFETA=700.007E+07;;;
+ MVST=800.008E+07
+ MXI=900.009E+07
+)

.model _3_PJF_PARKERSKELLERN pjf (level=2
+ VBI=000.000E+07;;;
+ AF=100.001E+07
+ BETA=200.002E+07
+ CDS=300.003E+07
+ CGD=400.004E+07
+ CGS=500.005E+07
+ DELTA=600.006E+07
+ HFETA=700.007E+07;;;
+ MVST=800.008E+07
+ MXI=900.009E+07
+)

.model _4_NMF_STATZ nmf (level=1
+ VTO=000.000E+07
+ ALPHA=100.001E+07
+ BETA=200.002E+07
+ LAMBDA=300.003E+07
+ B=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ CGS=700.007E+07
+ CGD=800.008E+07
+ PB=900.009E+07
+)

.model _5_PMF_STATZ pmf (level=1
+ VTO=000.000E+07
+ ALPHA=100.001E+07
+ BETA=200.002E+07
+ LAMBDA=300.003E+07
+ B=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ CGS=700.007E+07
+ CGD=800.008E+07
+ PB=900.009E+07
+)

* TODO: Ngspice User's Manual shows model line for MESFETs with level=4 - investigate that.
.model _6_NMF_YTTERDAL nmf (level=2
+ VTO=000.000E+07
+ LAMBDA=100.001E+07
+ LAMBDAHF=200.002E+07
+ BETA=300.003E+07
+ VS=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ RG=700.007E+07
+ RI=800.008E+07
+ RF=900.009E+07
+)

.model _7_PMF_YTTERDAL pmf (level=2
+ VTO=000.000E+07
+ LAMBDA=100.001E+07
+ LAMBDAHF=200.002E+07
+ BETA=300.003E+07
+ VS=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ RG=700.007E+07
+ RI=800.008E+07
+ RF=900.009E+07
+)

.model _8_NMF_HFET1 nmf (level=5
+ VTO=000.000E+07
+ LAMBDA=100.001E+07
+ RD=200.002E+07
+ RS=300.003E+07
+ RG=400.004E+07
+ RDI=500.005E+07
+ RSI=600.006E+07
+ RGS=700.007E+07
+ RGD=800.008E+07;;;
+ ETA=900.009E+07
+)

.model _9_PMF_HFET1 pmf (level=5
+ VTO=000.000E+07
+ LAMBDA=100.001E+07
+ RD=200.002E+07
+ RS=300.003E+07
+ RG=400.004E+07
+ RDI=500.005E+07
+ RSI=600.006E+07
+ RGS=700.007E+07
+ RGD=800.008E+07;;;
+ ETA=900.009E+07
+)

.model _10_NMF_HFET2 nmf (level=6
+ VS=000.000E+07;;;
+ GGR=100.001E+07
+ JS=200.002E+07;;;
+ DEL=300.003E+07
+ DELTA=400.004E+07
+ DELTAD=500.005E+07
+ DI=600.006E+07
+ EPSI=700.007E+07
+ ETA=800.008E+07
+ ETA1=900.009E+07
+)

.model _11_PMF_HFET2 pmf (level=6
+ VS=000.000E+07;;;
+ GGR=100.001E+07
+ JS=200.002E+07;;;
+ DEL=300.003E+07
+ DELTA=400.004E+07
+ DELTAD=500.005E+07
+ DI=600.006E+07
+ EPSI=700.007E+07
+ ETA=800.008E+07
+ ETA1=900.009E+07
+)

.model _12_NMOS_VD VDMOS NCHAN
*type, Not really a parameter.
+ vto         = 000.000E+07
*vth0, Alias.
+ kp          = 100.001E+07
+ phi         = 200.002E+07
+ lambda      = 300.003E+07
+ theta       = 400.004E+07
+ rd          = 500.005E+07
+ rs          = 600.006E+07
+ rg          = 700.007E+07
+ tnom        = 800.008E+07
+ kf          = 900.009E+07
+ af          = 000.000E+07
*vdmosn, Not really a parameter.
*vdmosp, Not really a parameter.
*vdmos, Not really a parameter.
+ rq          = 100.001E+07
+ vq          = 200.002E+07
+ mtriode     = 300.003E+07
+ tcvth       = 400.004E+07
*vtotc, Alias.
+ mu          = 500.005E+07
*bex, Alias.
+ texp0       = 600.006E+07
+ texp1       = 700.007E+07
+ trd1        = 800.008E+07
+ trd2        = 900.009E+07
+ trg1        = 000.000E+07
+ trg2        = 100.001E+07
+ trs1        = 200.002E+07
+ trs2        = 300.003E+07
+ trb1        = 400.004E+07
+ trb2        = 500.005E+07
+ subshift    = 600.006E+07
+ ksubthres   = 700.007E+07
+ tksubthres1 = 800.008E+07
+ tksubthres2 = 900.009E+07
+ bv          = 000.000E+07
+ ibv         = 100.001E+07
+ nbv         = 200.002E+07
+ rds         = 300.003E+07
+ rb          = 400.004E+07
+ n           = 500.005E+07
+ tt          = 600.006E+07
+ eg          = 700.007E+07
+ xti         = 800.008E+07
+ is          = 900.009E+07
+ vj          = 000.000E+07
+ cjo         = 100.001E+07
+ m           = 200.002E+07
+ fc          = 300.003E+07
+ cgdmin      = 400.004E+07
+ cgdmax      = 500.005E+07
+ a           = 600.006E+07
+ cgs         = 700.007E+07
+ rthjc       = 800.008E+07
+ rthca       = 900.009E+07
+ cthj        = 000.000E+07
+ vgs_max     = 100.001E+07
+ vgd_max     = 200.002E+07
+ vds_max     = 300.003E+07
+ vgsr_max    = 400.004E+07
+ vgdr_max    = 500.005E+07
+ pd_max      = 600.006E+07
+ id_max      = 700.007E+07
+ idr_max     = 800.008E+07
+ te_max      = 900.009E+07
+ rth_ext     = 000.000E+07
+ derating    = 100.001E+07 

.model _13_PMOS_VD VDMOS PCHAN
*type, Not really a parameter.
+ vto         = 000.000E+07
*vth0, Alias.
+ kp          = 100.001E+07
+ phi         = 200.002E+07
+ lambda      = 300.003E+07
+ theta       = 400.004E+07
+ rd          = 500.005E+07
+ rs          = 600.006E+07
+ rg          = 700.007E+07
+ tnom        = 800.008E+07
+ kf          = 900.009E+07
+ af          = 000.000E+07
*vdmosn, Not really a parameter.
*vdmosp, Not really a parameter.
*vdmos, Not really a parameter.
+ rq          = 100.001E+07
+ vq          = 200.002E+07
+ mtriode     = 300.003E+07
+ tcvth       = 400.004E+07
*vtotc, Alias.
+ mu          = 500.005E+07
*bex, Alias.
+ texp0       = 600.006E+07
+ texp1       = 700.007E+07
+ trd1        = 800.008E+07
+ trd2        = 900.009E+07
+ trg1        = 000.000E+07
+ trg2        = 100.001E+07
+ trs1        = 200.002E+07
+ trs2        = 300.003E+07
+ trb1        = 400.004E+07
+ trb2        = 500.005E+07
+ subshift    = 600.006E+07
+ ksubthres   = 700.007E+07
+ tksubthres1 = 800.008E+07
+ tksubthres2 = 900.009E+07
+ bv          = 000.000E+07
+ ibv         = 100.001E+07
+ nbv         = 200.002E+07
+ rds         = 300.003E+07
+ rb          = 400.004E+07
+ n           = 500.005E+07
+ tt          = 600.006E+07
+ eg          = 700.007E+07
+ xti         = 800.008E+07
+ is          = 900.009E+07
+ vj          = 000.000E+07
+ cjo         = 100.001E+07
+ m           = 200.002E+07
+ fc          = 300.003E+07
+ cgdmin      = 400.004E+07
+ cgdmax      = 500.005E+07
+ a           = 600.006E+07
+ cgs         = 700.007E+07
+ rthjc       = 800.008E+07
+ rthca       = 900.009E+07
+ cthj        = 000.000E+07
+ vgs_max     = 100.001E+07
+ vgd_max     = 200.002E+07
+ vds_max     = 300.003E+07
+ vgsr_max    = 400.004E+07
+ vgdr_max    = 500.005E+07
+ pd_max      = 600.006E+07
+ id_max      = 700.007E+07
+ idr_max     = 800.008E+07
+ te_max      = 900.009E+07
+ rth_ext     = 000.000E+07
+ derating    = 100.001E+07 

.model _14_NMOS_MOS1 nmos (level=1
+ VTO=000.000E+07
+ KP=100.001E+07
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ LAMBDA=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _15_PMOS_MOS1 pmos (level=1
+ VTO=000.000E+07
+ KP=100.001E+07
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ LAMBDA=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _16_NMOS_MOS2 nmos (level=2
+ VTO=000.000E+07
+ KP=100.001E+07
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ LAMBDA=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _17_PMOS_MOS2 pmos (level=2
+ VTO=000.000E+07
+ KP=100.001E+07 ; Does not exist in MOS3 and MOS6
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ LAMBDA=400.004E+07 ; Does not exist in MOS3
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _18_NMOS_MOS3 nmos (level=3
+ VTO=000.000E+07
+ THETA=100.001E+07 ; MOS3 and MOS9-only
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ ETA=400.004E+07 ; MOS3 and MOS9-only
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _19_PMOS_MOS3 pmos (level=3
+ VTO=000.000E+07
+ THETA=100.001E+07 ; MOS3 and MOS9-only
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ ETA=400.004E+07 ; MOS3 and MOS9-only
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _20_NMOS_BSIM1 nmos (level=4
+ VFB=000.000E+07
+ LVFB=100.001E+07
+ WVFB=200.002E+07
+ PHI=300.003E+07
+ LPHI=400.004E+07
+ WPHI=500.005E+07
+ K1=600.006E+07
+ LK1=700.007E+07
+ WK1=800.008E+07
+ K2=900.009E+07
+)

.model _21_PMOS_BSIM1 pmos (level=4
+ VFB=000.000E+07
+ LVFB=100.001E+07
+ WVFB=200.002E+07
+ PHI=300.003E+07
+ LPHI=400.004E+07
+ WPHI=500.005E+07
+ K1=600.006E+07
+ LK1=700.007E+07
+ WK1=800.008E+07
+ K2=900.009E+07
+)

.model _22_NMOS_BSIM2 nmos (level=5
+ BIB=000.000E+07
+ LBIB=100.001E+07
+ WBIB=200.002E+07
+ VGHIGH=300.003E+07
+ LVGHIGH=400.004E+07
+ WVGHIGH=500.005E+07;;;
+ WAIB=600.006E+07
+ BI0=700.007E+07
+ LBI0=800.008E+07
+ WBI0=900.009E+07
+)

.model _23_PMOS_BSIM2 pmos (level=5
+ BIB=000.000E+07
+ LBIB=100.001E+07
+ WBIB=200.002E+07
+ VGHIGH=300.003E+07
+ LVGHIGH=400.004E+07
+ WVGHIGH=500.005E+07;;;
+ WAIB=600.006E+07
+ BI0=700.007E+07
+ LBI0=800.008E+07
+ WBI0=900.009E+07
+)

.model _24_NMOS_MOS6 nmos (level=6
+ VTO=000.000E+07
+ NVTH=100.001E+07 ; MOS6-only
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ LAMBDA=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _25_PMOS_MOS6 pmos (level=6
+ VTO=000.000E+07
+ NVTH=100.001E+07 ; MOS6-only
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ LAMBDA=400.004E+07
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _26_NMOS_BSIM3 nmos (level=8
+ TOX=000.000E+07
+ TOXM=100.001E+07
+ CDSC=200.002E+07
+ CDSCB=300.003E+07
+ CDSCD=400.004E+07
+ CIT=500.005E+07
+ NFACTOR=600.006E+07
+ XJ=700.007E+07
+ VSAT=800.008E+07
+ AT=900.009E+07
+)

.model _27_PMOS_BSIM3 pmos (level=8
+ TOX=000.000E+07
+ TOXM=100.001E+07
+ CDSC=200.002E+07
+ CDSCB=300.003E+07
+ CDSCD=400.004E+07
+ CIT=500.005E+07
+ NFACTOR=600.006E+07
+ XJ=700.007E+07
+ VSAT=800.008E+07
+ AT=900.009E+07
+)

.model _28_NMOS_MOS9 nmos (level=9
+ VTO=000.000E+07
+ THETA=100.001E+07 ; MOS3 and MOS9-only
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ ETA=400.004E+07 ; MOS3 and MOS9-only
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _29_PMOS_MOS9 pmos (level=9
+ VTO=000.000E+07
+ THETA=100.001E+07 ; MOS3 and MOS9-only
+ GAMMA=200.002E+07
+ PHI=300.003E+07
+ ETA=400.004E+07 ; MOS3 and MOS9-only
+ RD=500.005E+07
+ RS=600.006E+07
+ CBD=700.007E+07
+ CBS=800.008E+07
+ IS=900.009E+07
+)

.model _30_NMOS_B4SOI nmos (level=10
+ TOX=000.000E+07
+ TOXP=100.001E+07
+ TOXM=200.002E+07
+ DTOXCV=300.003E+07
+ CDSC=400.004E+07
+ CDSCB=500.005E+07
+ CDSCD=600.006E+07
+ CIT=700.007E+07
+ NFACTOR=800.008E+07
+ VSAT=900.009E+07
+)

.model _31_PMOS_B4SOI pmos (level=10
+ TOX=000.000E+07
+ TOXP=100.001E+07
+ TOXM=200.002E+07
+ DTOXCV=300.003E+07
+ CDSC=400.004E+07
+ CDSCB=500.005E+07
+ CDSCD=600.006E+07
+ CIT=700.007E+07
+ NFACTOR=800.008E+07
+ VSAT=900.009E+07
+)

.model _32_NMOS_BSIM4 nmos (level=14
+ RBPS0=000.000E+07
+ RBPSL=100.001E+07
+ RBPSW=200.002E+07
+ RBPSNF=300.003E+07
+ RBPD0=400.004E+07
+ RBPDL=500.005E+07
+ RBPDW=600.006E+07
+ RBPDNF=700.007E+07
+ RBPBX0=800.008E+07
+ RBPBXL=900.009E+07
+)

.model _33_PMOS_BSIM4 pmos (level=14
+ RBPS0=000.000E+07
+ RBPSL=100.001E+07
+ RBPSW=200.002E+07
+ RBPSNF=300.003E+07
+ RBPD0=400.004E+07
+ RBPDL=500.005E+07
+ RBPDW=600.006E+07
+ RBPDNF=700.007E+07
+ RBPBX0=800.008E+07
+ RBPBXL=900.009E+07
+)

.model _34_NMOS_B3SOIFD nmos (level=55
+ TOX=000.000E+07
+ CDSC=100.001E+07
+ CDSCB=200.002E+07
+ CDSCD=300.003E+07
+ CIT=400.004E+07
+ NFACTOR=500.005E+07
+ VSAT=600.006E+07
+ AT=700.007E+07
+ A0=800.008E+07
+ AGS=900.009E+07
+)

.model _35_PMOS_B3SOIFD pmos (level=55
+ TOX=000.000E+07
+ CDSC=100.001E+07
+ CDSCB=200.002E+07
+ CDSCD=300.003E+07
+ CIT=400.004E+07
+ NFACTOR=500.005E+07
+ VSAT=600.006E+07
+ AT=700.007E+07
+ A0=800.008E+07
+ AGS=900.009E+07
+)

.model _36_NMOS_B3SOIDD nmos (level=56
+ TOX=000.000E+07
+ CDSC=100.001E+07
+ CDSCB=200.002E+07
+ CDSCD=300.003E+07
+ CIT=400.004E+07
+ NFACTOR=500.005E+07
+ VSAT=600.006E+07
+ AT=700.007E+07
+ A0=800.008E+07
+ AGS=900.009E+07
+)

.model _37_PMOS_B3SOIDD pmos (level=56
+ TOX=000.000E+07
+ CDSC=100.001E+07
+ CDSCB=200.002E+07
+ CDSCD=300.003E+07
+ CIT=400.004E+07
+ NFACTOR=500.005E+07
+ VSAT=600.006E+07
+ AT=700.007E+07
+ A0=800.008E+07
+ AGS=900.009E+07
+)

.model _38_NMOS_B3SOIPD nmos (level=57
+ TOX=000.000E+07
+ CDSC=100.001E+07
+ CDSCB=200.002E+07
+ CDSCD=300.003E+07
+ CIT=400.004E+07
+ NFACTOR=500.005E+07
+ VSAT=600.006E+07
+ AT=700.007E+07
+ A0=800.008E+07
+ AGS=900.009E+07
+)

.model _39_PMOS_B3SOIPD pmos (level=57
+ TOX=000.000E+07
+ CDSC=100.001E+07
+ CDSCB=200.002E+07
+ CDSCD=300.003E+07
+ CIT=400.004E+07
+ NFACTOR=500.005E+07
+ VSAT=600.006E+07
+ AT=700.007E+07
+ A0=800.008E+07
+ AGS=900.009E+07
+)

.model _40_NMOS_HISIM2 nmos (level=68
+ DEPMUE0=000.000E+07
+ DEPMUE0L=100.001E+07
+ DEPMUE0LP=200.002E+07
+ DEPMUE1=300.003E+07
+ DEPMUE1L=400.004E+07
+ DEPMUE1LP=500.005E+07
+ DEPMUEBACK0=600.006E+07
+ DEPMUEBACK0L=700.007E+07
+ DEPMUEBACK0LP=800.008E+07
+ DEPMUEBACK1=900.009E+07
+)

.model _41_PMOS_HISIM2 pmos (level=68
+ DEPMUE0=000.000E+07
+ DEPMUE0L=100.001E+07
+ DEPMUE0LP=200.002E+07
+ DEPMUE1=300.003E+07
+ DEPMUE1L=400.004E+07
+ DEPMUE1LP=500.005E+07
+ DEPMUEBACK0=600.006E+07
+ DEPMUEBACK0L=700.007E+07
+ DEPMUEBACK0LP=800.008E+07
+ DEPMUEBACK1=900.009E+07
+)

.model _42_NMOS_HISIMHV1 nmos (level=73 version=1.2.4
+ PRD=000.000E+07
+ PRD22=100.001E+07
+ PRD23=200.002E+07
+ PRD24=300.003E+07
+ PRDICT1=400.004E+07
+ PRDOV13=500.005E+07
+ PRDSLP1=600.006E+07
+ PRDVB=700.007E+07
+ PRDVD=800.008E+07
+ PRDVG11=900.009E+07
+)

.model _43_PMOS_HISIMHV1 pmos (level=73 version=1.2.4
+ PRD=000.000E+07
+ PRD22=100.001E+07
+ PRD23=200.002E+07
+ PRD24=300.003E+07
+ PRDICT1=400.004E+07
+ PRDOV13=500.005E+07
+ PRDSLP1=600.006E+07
+ PRDVB=700.007E+07
+ PRDVD=800.008E+07
+ PRDVG11=900.009E+07
+)

.model _44_NMOS_HISIMHV2 nmos (level=73 version=2.2.0
+ PJS0D=000.000E+07
+ PJS0SWD=100.001E+07
+ PNJD=200.002E+07
+ PCISBKD=300.003E+07
+ PVDIFFJD=400.004E+07
+ PJS0S=500.005E+07
+ PJS0SWS=600.006E+07;;;
+ PRS=700.007E+07
+ PRTH0=800.008E+07
+ PVOVER=900.009E+07
+)

.model _45_PMOS_HISIMHV2 pmos (level=73 version=2.2.0
+ PJS0D=000.000E+07
+ PJS0SWD=100.001E+07
+ PNJD=200.002E+07
+ PCISBKD=300.003E+07
+ PVDIFFJD=400.004E+07
+ PJS0S=500.005E+07
+ PJS0SWS=600.006E+07;;;
+ PRS=700.007E+07
+ PRTH0=800.008E+07
+ PVOVER=900.009E+07
+)
