��ࡱ�                >  ��	                               ����        ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������            	   ����   
   ����                  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������R o o t   E n t r y                                               ��������                               p�� |�   �      C a c h e                                                        ������������                                    !   
       C e l l s                                                              ����                    p�� |�p�� |�            P a r t s                                                        ������������                    p�� |�p�� |�            V i e w s                                                               ����                    p�� |�p�� |�            L i b r a r y                                                    ������������                                    	   �      S y m b o l s                                                                                 p�� |�p�� |�            G r a p h i c s                                                  ��������                       p�� |�p�� |�            P a c k a g e s                                                                               p�� |�p�� |�            E x p o r t B l o c k s                                          ������������                    p�� |�p�� |�            C e l l s   D i r e c t o r y                                     	      ����                                       &       P a r t s   D i r e c t o r y                                     ������������                                       U       V i e w s   D i r e c t o r y                                      
      ����                                              N e t B u n d l e M a p D a t a                                 " ������������                                              S y m b o l s   D i r e c t o r y                               $       ����                                              G r a p h i c s   D i r e c t o r y                             &  ������������                                              P a c k a g e s   D i r e c t o r y                             &       ����                                       &       E x p o r t B l o c k s   D i r e c t o r y                     .  ������������                                               O P A 1 6 4 x                                                    ������������                                    "   	      $ T y p e s $                                                    ������������                                    ����        ������������������������   ��������
                                                                      ��������#   $   %   &   '   (   )   *   +   ,   -   .   /   0   1   2   3   4   5   6   7   8   9   :   ;   <   =   >   ?   @   A   B   ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������P#�b           IN-        ����   !               VP#�b  OPA164x  `�8N|� 
�8N|��   Amp6T_TI  бt�V�@4xP#�b    Amp6B_TI  ��7�V� P��V��  Amp9_TI  vo\���P#�b  �  Amp7_TI  0M��[��@��[��  Amp5_TI   �kJZ�0�   �� 	 InAmp8_TI   %��U����U��  2  5  3  4  P#�b   OPA2333P  ���)�� �[V+��                            P#�b  OPA164x.Normal  `�8N|� 
�8N|��  OPA164x.Convert  �`�8N|� 
�8N|�� mal   %��U����U��  Amp6B_TI.NormalP#�b  OPA164x  `�8N|� 
�8N|�� �U��  Amp6B_TI.NormalOrCAD Windows Library             �.H\P#�b    
 ����           �      "Arial �ei ����9� ��t�����           �      1Courier New l���cYt��              �     �  Arial �b          OPA333.Norma              �     � Arial �/              OiTH֌/����            �      Arial ng package..Amp5_TI       ����            �      Arial mp\CDN_SYMEDITOR_temp.olb ����           �     � Arial %+ %$ T y p e s $                                                    ������������                                    ����                                                                            ������������                                                                                                                    ������������                                                                                                                    ������������                                                - %V+ %V- %OUT @MODEL ����            �      Arial %+ %- %V+ %V- %OUT @MODEL ����            �      Arial %+ %- %V+ %V- %OUT @MODEL                                            1ST PART FIELD  2ND PART FIELD  3RD PART FIELD  4TH PART FIELD  5TH PART FIELD  6TH PART FIELD  7TH PART FIELD  PCB Footprint                                 d         d   d   0   0                                                                                                 Part Reference  Value  PSpiceTemplate * X^@REFDES %IN+ %IN- %VCC %VEE %OUT @MODEL   FLOAT  Error ) X^@REFDES %IN+ %IN- %VCC %VEE %OUT @MODEL # X^@REFDES %+ %- %V+ %V- %OUT @MODEL  Name 6 X^@REFDES %IN+ %IN- %RG+ %RG- %V+ %V- %OUT %REF @MODEL ' X^@REFDES %+ %- %V+ %V- %OUT %SD @MODEL ' X^@REFDES %+ %- %V+ %V- %OUT %EN @MODEL ( X^@REFDES %+ %- %V+ %V- %OUT %REF @MODEL C X^@REFDES %+ %- %V+ %V- %OUT %P1 %P2 %P3 %P4 %P1 %P2 %P3 %P4 @MODEL 3 X^@REFDES %+ %- %V+ %V- %OUT %P1 %P2 %P3 %P4 @MODEL 0 X^@REFDES %+ %- %V+ %V- %OUT+ %OUT- %VOCM @MODEL   �cYt��              �              l �b          OPA333.Norma              �     �  O       !              ����\9     OPA164x      OPA164x.Normal  OPA164x.Convert  �      e            0                     ��\9     OPA164x.Normal    0    ))                <             ��\9    ))        <          <          ��\9    ))                    <          ��\9    ))                             ��\9    ))           <      -           ��\9        < <  >                     ��\9     +     
   ����
   !           >                     ��\9     -     2   ����2   !           j                     ��\9     V+               !          '"       '       '����\9    	        0  j                     ��\9     V-    <      <   !          '"       '       '����\9    	     .   0  @                     ��\9     OUT <      F      !            '8       '!       '����\9            2 47 -5      + �� 0  '8       '!       '����\9            2 58 64      + =  0      OPA164X  U  OPA164x / �      f            1                     ��\9     OPA164x.Convert    0    ))        <          <          ��\9    ))                    <          ��\9    ))                <             ��\9    ))                             ��\9    ))           <      -           ��\9        < <  >                     ��\9     +     2   ����2   !           >                     ��\9     -     
   ����
   ! o     I   j                     ��\9     V+               !       e  '"       '       '����\9    	        0  j                     ��\9     V-    <      <   !          '"       '       '����\9    	   ! /   0  @                     ��\9     OUT <      F      !       L    '8       '!       '����\9            2 47 -5      + �� 0  '8       '!       '����\9            2 58 64      + =  0      OPA164x  U  OPA164x / {       !                ��\9     OPA164x     U         <                ����\9        OPA164x   1  2  5  3  4                                                                                                                                                                                                                                                                                                                                                                                        