* EESchema Netlist Version 1.1 (Spice format) creation date: 14/07/2010 14:49:50


R12  VOUT N-000010 22K
R11  +12V N-000010 100
L1  N-000010 VOUT 100mH
R10  N-000009 N-000004 220
C3  N-000009 0 10uF
C2  N-000008 0 1nF
R8  N-000004 0 2.2K
Q3  VOUT N-000008 N-000004 N-000004 Q2N2222
V2  N-000003 0 AC 0.1
C1  VIN N-000003 1UF
V1  +12V 0 DC 12V
R2  VIN 0 10K
R6  +12V VIN 22K
R5  +12V N-000006 22K
R1  N-000006 0 10K
R7  N-000005 0 470
R4  +12V N-000008 1K
R3  +12V N-000007 1K
Q2  N-000008 N-000006 N-000005 N-000005 Q2N2222
Q1  N-000007 VIN N-000005 N-000005 Q2N2222

.model Q2N2222 npn (bf=200)
.print tran v(nodes)
.print dc v(nodes)
.tran 10 10000 10 > x.txt
.save all

.end
