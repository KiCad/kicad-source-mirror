*
* bjts.lib.spice
* 

* All parameter values are made up and physically nonsensical.
* Commented out some parameters to avoid making test code overly long.


* VBIC.

.model _0_NPN_VBIC NPN( level=4
+ rcx             = 000.000E+07
+ rci             = 100.001E+07
+ vo              = 200.002E+07
+ gamm            = 300.003E+07
+ hrcf            = 400.004E+07
+ rbx             = 500.005E+07
+ rbi             = 600.006E+07
+ re              = 700.007E+07
+ rs              = 800.008E+07
+ rbp             = 900.009E+07
+ is              = 000.000E+07
+ nf              = 100.001E+07
+ nr              = 200.002E+07
+ fc              = 300.003E+07
+ cbeo            = 400.004E+07
+ cje             = 500.005E+07
+ pe              = 600.006E+07
+ me              = 700.007E+07
+ aje             = 800.008E+07
+ cbco            = 900.009E+07
+ cjc             = 000.000E+07
+ qco             = 100.001E+07
+ cjep            = 200.002E+07
+ pc              = 300.003E+07
+ mc              = 400.004E+07
+ ajc             = 500.005E+07
+ cjcp            = 600.006E+07
+ ps              = 700.007E+07
+ ms              = 800.008E+07
+ ajs             = 900.009E+07
+ ibei            = 000.000E+07
+ wbe             = 100.001E+07
+ nei             = 200.002E+07
+ iben            = 300.003E+07
+ nen             = 400.004E+07
+ ibci            = 500.005E+07
+ nci             = 600.006E+07
+ ibcn            = 700.007E+07
+ ncn             = 800.008E+07
+ avc1            = 900.009E+07
+ avc2            = 000.000E+07
+ isp             = 100.001E+07
+ wsp             = 200.002E+07
+ nfp             = 300.003E+07
+ ibeip           = 400.004E+07
+ ibenp           = 500.005E+07
+ ibcip           = 600.006E+07
+ ncip            = 700.007E+07
+ ibcnp           = 800.008E+07
+ ncnp            = 900.009E+07
+ vef             = 000.000E+07
+ ver             = 100.001E+07
+ ikf             = 200.002E+07
+ ikr             = 300.003E+07
+ ikp             = 400.004E+07
+ tf              = 500.005E+07
+ qtf             = 600.006E+07
+ xtf             = 700.007E+07
+ vtf             = 800.008E+07
+ itf             = 900.009E+07
+ tr              = 000.000E+07
+ td              = 100.001E+07
+ kfn             = 200.002E+07
+ afn             = 300.003E+07
+ bfn             = 400.004E+07
+ xre             = 500.005E+07
+ xrb             = 600.006E+07
+ xrbi            = 700.007E+07
+ xrc             = 800.008E+07
+ xrci            = 900.009E+07
+ xrs             = 000.000E+07
+ xvo             = 100.001E+07
+ ea              = 200.002E+07
+ eaie            = 300.003E+07
+ eaic            = 400.004E+07
+ eais            = 500.005E+07
+ eane            = 600.006E+07
+ eanc            = 700.007E+07
+ eans            = 800.008E+07
+ xis             = 900.009E+07
+ xii             = 000.000E+07
+ xin             = 100.001E+07
+ tnf             = 200.002E+07
+ tavc            = 300.003E+07
+ rth             = 400.004E+07
+ cth             = 500.005E+07
+ vrt             = 600.006E+07
+ art             = 700.007E+07
+ ccso            = 800.008E+07
+ qbm             = 900.009E+07
+ nkf             = 000.000E+07
+ xikf            = 100.001E+07
+ xrcx            = 200.002E+07
+ xrbx            = 300.003E+07
+ xrbp            = 400.004E+07
+ isrr            = 500.005E+07
+ xisr            = 600.006E+07
+ dear            = 700.007E+07
+ eap             = 800.008E+07
+ vbbe            = 900.009E+07
+ nbbe            = 000.000E+07
+ ibbe            = 100.001E+07
+ tvbbe1          = 200.002E+07
+ tvbbe2          = 300.003E+07
+ tnbbe           = 400.004E+07
+ ebbe            = 500.005E+07
+ dtemp           = 600.006E+07
+ vers            = 700.007E+07
+ vref            = 800.008E+07
+ vbe_max         = 900.009E+07
+ vbc_max         = 000.000E+07
+ vce_max         = 100.001E+07
+)

.model _1_PNP_VBIC PNP( level=4.0
+ rcx             = 000.000E+07
+ rci             = 100.001E+07
+ vo              = 200.002E+07
+ gamm            = 300.003E+07
+ hrcf            = 400.004E+07
+ rbx             = 500.005E+07
+ rbi             = 600.006E+07
+ re              = 700.007E+07
+ rs              = 800.008E+07
+ rbp             = 900.009E+07
+ is              = 000.000E+07
+ nf              = 100.001E+07
+ nr              = 200.002E+07
+ fc              = 300.003E+07
+ cbeo            = 400.004E+07
+ cje             = 500.005E+07
+ pe              = 600.006E+07
+ me              = 700.007E+07
+ aje             = 800.008E+07
+ cbco            = 900.009E+07
+ cjc             = 000.000E+07
+ qco             = 100.001E+07
+ cjep            = 200.002E+07
+ pc              = 300.003E+07
+ mc              = 400.004E+07
+ ajc             = 500.005E+07
+ cjcp            = 600.006E+07
+ ps              = 700.007E+07
+ ms              = 800.008E+07
+ ajs             = 900.009E+07
+ ibei            = 000.000E+07
+ wbe             = 100.001E+07
+ nei             = 200.002E+07
+ iben            = 300.003E+07
+ nen             = 400.004E+07
+ ibci            = 500.005E+07
+ nci             = 600.006E+07
+ ibcn            = 700.007E+07
+ ncn             = 800.008E+07
+ avc1            = 900.009E+07
+ avc2            = 000.000E+07
+ isp             = 100.001E+07
+ wsp             = 200.002E+07
+ nfp             = 300.003E+07
+ ibeip           = 400.004E+07
+ ibenp           = 500.005E+07
+ ibcip           = 600.006E+07
+ ncip            = 700.007E+07
+ ibcnp           = 800.008E+07
+ ncnp            = 900.009E+07
+ vef             = 000.000E+07
+ ver             = 100.001E+07
+ ikf             = 200.002E+07
+ ikr             = 300.003E+07
+ ikp             = 400.004E+07
+ tf              = 500.005E+07
+ qtf             = 600.006E+07
+ xtf             = 700.007E+07
+ vtf             = 800.008E+07
+ itf             = 900.009E+07
+ tr              = 000.000E+07
+ td              = 100.001E+07
+ kfn             = 200.002E+07
+ afn             = 300.003E+07
+ bfn             = 400.004E+07
+ xre             = 500.005E+07
+ xrb             = 600.006E+07
+ xrbi            = 700.007E+07
+ xrc             = 800.008E+07
+ xrci            = 900.009E+07
+ xrs             = 000.000E+07
+ xvo             = 100.001E+07
+ ea              = 200.002E+07
+ eaie            = 300.003E+07
+ eaic            = 400.004E+07
+ eais            = 500.005E+07
+ eane            = 600.006E+07
+ eanc            = 700.007E+07
+ eans            = 800.008E+07
+ xis             = 900.009E+07
+ xii             = 000.000E+07
+ xin             = 100.001E+07
+ tnf             = 200.002E+07
+ tavc            = 300.003E+07
+ rth             = 400.004E+07
+ cth             = 500.005E+07
+ vrt             = 600.006E+07
+ art             = 700.007E+07
+ ccso            = 800.008E+07
+ qbm             = 900.009E+07
+ nkf             = 000.000E+07
+ xikf            = 100.001E+07
+ xrcx            = 200.002E+07
+ xrbx            = 300.003E+07
+ xrbp            = 400.004E+07
+ isrr            = 500.005E+07
+ xisr            = 600.006E+07
+ dear            = 700.007E+07
+ eap             = 800.008E+07
+ vbbe            = 900.009E+07
+ nbbe            = 000.000E+07
+ ibbe            = 100.001E+07
+ tvbbe1          = 200.002E+07
+ tvbbe2          = 300.003E+07
+ tnbbe           = 400.004E+07
+ ebbe            = 500.005E+07
+ dtemp           = 600.006E+07
+ vers            = 700.007E+07
+ vref            = 800.008E+07
+ vbe_max         = 900.009E+07
+ vbc_max         = 000.000E+07
+ vce_max         = 100.001E+07
+)


* SPICE Gummel-Poon.

*
.MODEL _2_NPN_GUMMELPOON NPN(  
+     IS   = 000.000E+07
+     NF   = 100.001E+07
+     ISE  = 200.002E+07
+     NE   = 300.003E+07
+     BF   = 400.004E+07
+     IKF  = 500.005E+07
+     VAF  = 600.006E+07
+     NR   = 700.007E+07
+     ISC  = 800.008E+07
+     NC   = 900.009E+07
+     BR   = 000.000E+07
+     IKR  = 100.001E+07
+     VAR  = 200.002E+07
+     RB   = 300.003E+07
+     IRB  = 400.004E+07
+     RBM  = 500.005E+07
+     RE   = 600.006E+07
+     RC   = 700.007E+07
+     XTB  = 800.008E+07
+     EG   = 900.009E+07
+     XTI  = 000.000E+07
+     CJE  = 100.001E+07
+     VJE  = 200.002E+07
+     MJE  = 300.003E+07
+     TF   = 400.004E+07
+     XTF  = 500.005E+07
+     VTF  = 600.006E+07
+     ITF  = 700.007E+07
+     PTF  = 800.008E+07
+     CJC  = 900.009E+07
+     VJC  = 000.000E+07
+     MJC  = 100.001E+07
+     XCJC = 200.002E+07
+     TR   = 300.003E+07
+     CJS  = 400.004E+07
+     VJS  = 500.005E+07
+     MJS  = 600.006E+07
+     FC   = 700.007E+07
+)


*
.MODEL _3_PNP_GUMMELPOON PNP( level = 1. ; Decimal separator must be accepted too.
+     IS   = 000.000E+07
+     NF   = 100.001E+07
+     ISE  = 200.002E+07
+     NE   = 300.003E+07
+     BF   = 400.004E+07
+     IKF  = 500.005E+07
+     VAF  = 600.006E+07
+     NR   = 700.007E+07
+     ISC  = 800.008E+07
+     NC   = 900.009E+07
+     BR   = 000.000E+07
+     IKR  = 100.001E+07
+     VAR  = 200.002E+07
+     RB   = 300.003E+07
+     IRB  = 400.004E+07
+     RBM  = 500.005E+07
+     RE   = 600.006E+07
+     RC   = 700.007E+07
+     XTB  = 800.008E+07
+     EG   = 900.009E+07
+     XTI  = 000.000E+07
+     CJE  = 100.001E+07
+     VJE  = 200.002E+07
+     MJE  = 300.003E+07
+     TF   = 400.004E+07
+     XTF  = 500.005E+07
+     VTF  = 600.006E+07
+     ITF  = 700.007E+07
+     PTF  = 800.008E+07
+     CJC  = 900.009E+07
+     VJC  = 000.000E+07
+     MJC  = 100.001E+07
+     XCJC = 200.002E+07
+     TR   = 300.003E+07
+     CJS  = 400.004E+07
+     VJS  = 500.005E+07
+     MJS  = 600.006E+07
+     FC   = 700.007E+07
+)


* HICUM/L2.

.model _4_NPN_HICUML2 NPN( level=8.00
+ c10             = 000.000E+07
+ qp0             = 100.001E+07
+ ich             = 200.002E+07
+ hf0             = 300.003E+07
+ hfe             = 400.004E+07
+ hfc             = 500.005E+07
+ hjei            = 600.006E+07
+ ahjei           = 700.007E+07
+ rhjei           = 800.008E+07
+ hjci            = 900.009E+07
+ ibeis           = 000.000E+07
+ mbei            = 100.001E+07
+ ireis           = 200.002E+07
+ mrei            = 300.003E+07
+ ibeps           = 400.004E+07
+ mbep            = 500.005E+07
+ ireps           = 600.006E+07
+ mrep            = 700.007E+07
+ mcf             = 800.008E+07
+ tbhrec          = 900.009E+07
+ ibcis           = 000.000E+07
+ mbci            = 100.001E+07
+ ibcxs           = 200.002E+07
+ mbcx            = 300.003E+07
+ ibets           = 400.004E+07
+ abet            = 500.005E+07
+ tunode          = 6
+ favl            = 700.007E+07
+ qavl            = 800.008E+07
+ kavl            = 900.009E+07
+ alfav           = 000.000E+07
+ alqav           = 100.001E+07
+ alkav           = 200.002E+07
+ rbi0            = 300.003E+07
+ rbx             = 400.004E+07
+ fgeo            = 500.005E+07
+ fdqr0           = 600.006E+07
+ fcrbi           = 700.007E+07
+ fqi             = 800.008E+07
+ re              = 900.009E+07
+ rcx             = 000.000E+07
+ itss            = 100.001E+07
+ msf             = 200.002E+07
+ iscs            = 300.003E+07
+ msc             = 400.004E+07
+ tsf             = 500.005E+07
+ rsu             = 600.006E+07
+ csu             = 700.007E+07
+ cjei0           = 800.008E+07
+ vdei            = 900.009E+07
+ zei             = 000.000E+07
+ ajei            = 100.001E+07
*aljei
+ cjep0           = 200.002E+07
+ vdep            = 300.003E+07
+ zep             = 400.004E+07
+ ajep            = 500.005E+07
*aljep
+ cjci0           = 600.006E+07
+ vdci            = 700.007E+07
+ zci             = 800.008E+07
+ vptci           = 900.009E+07
+ cjcx0           = 000.000E+07
+ vdcx            = 100.001E+07
+ zcx             = 200.002E+07
+ vptcx           = 300.003E+07
+ fbcpar          = 400.004E+07
*+ fbc
+ fbepar          = 500.005E+07
*+ fbe
+ cjs0            = 600.006E+07
+ vds             = 700.007E+07
+ zs              = 800.008E+07
+ vpts            = 900.009E+07
+ cscp0           = 000.000E+07
+ vdsp            = 100.001E+07
+ zsp             = 200.002E+07
+ vptsp           = 300.003E+07
+ t0              = 400.004E+07
+ dt0h            = 500.005E+07
+ tbvl            = 600.006E+07
+ tef0            = 700.007E+07
+ gtfe            = 800.008E+07
+ thcs            = 900.009E+07
+ ahc             = 000.000E+07
*alhc
+ fthc            = 100.001E+07
+ rci0            = 200.002E+07
+ vlim            = 300.003E+07
+ vces            = 400.004E+07
+ vpt             = 500.005E+07
+ aick            = 600.006E+07
+ delck           = 700.007E+07
+ tr              = 800.008E+07
+ vcbar           = 900.009E+07
+ icbar           = 000.000E+07
+ acbar           = 100.001E+07
+ cbepar          = 200.002E+07
*ceox
+ cbcpar          = 300.003E+07
*ccox
+ alqf            = 400.004E+07
+ alit            = 500.005E+07
+ flnqs           = 6
+ kf              = 700.007E+07
+ af              = 800.008E+07
+ cfbe            = 9
+ flcono          = 0
+ kfre            = 100.001E+07
+ afre            = 200.002E+07
+ latb            = 300.003E+07
+ latl            = 400.004E+07
+ vgb             = 500.005E+07
+ alt0            = 600.006E+07
+ kt0             = 700.007E+07
+ zetaci          = 800.008E+07
+ alvs            = 900.009E+07
+ alces           = 000.000E+07
+ zetarbi         = 100.001E+07
+ zetarbx         = 200.002E+07
+ zetarcx         = 300.003E+07
+ zetare          = 400.004E+07
+ zetacx          = 500.005E+07
+ vge             = 600.006E+07
+ vgc             = 700.007E+07
+ vgs             = 800.008E+07
+ f1vg            = 900.009E+07
+ f2vg            = 000.000E+07
+ zetact          = 100.001E+07
+ zetabet         = 200.002E+07
+ alb             = 300.003E+07
+ dvgbe           = 400.004E+07
+ zetahjei        = 500.005E+07
+ zetavgbe        = 600.006E+07
+ flsh            = 7
+ rth             = 800.008E+07
+ zetarth         = 900.009E+07
+ alrth           = 000.000E+07
+ cth             = 100.001E+07
+ flcomp          = 200.002E+07
+ vbe_max         = 300.003E+07
+ vbc_max         = 400.004E+07
+ vce_max         = 500.005E+07
+)

.model _5_PNP_HICUML2 PNP( level=8
+ c10             = 000.000E+07
+ qp0             = 100.001E+07
+ ich             = 200.002E+07
+ hf0             = 300.003E+07
+ hfe             = 400.004E+07
+ hfc             = 500.005E+07
+ hjei            = 600.006E+07
+ ahjei           = 700.007E+07
+ rhjei           = 800.008E+07
+ hjci            = 900.009E+07
+ ibeis           = 000.000E+07
+ mbei            = 100.001E+07
+ ireis           = 200.002E+07
+ mrei            = 300.003E+07
+ ibeps           = 400.004E+07
+ mbep            = 500.005E+07
+ ireps           = 600.006E+07
+ mrep            = 700.007E+07
+ mcf             = 800.008E+07
+ tbhrec          = 900.009E+07
+ ibcis           = 000.000E+07
+ mbci            = 100.001E+07
+ ibcxs           = 200.002E+07
+ mbcx            = 300.003E+07
+ ibets           = 400.004E+07
+ abet            = 500.005E+07
+ tunode          = 6
+ favl            = 700.007E+07
+ qavl            = 800.008E+07
+ kavl            = 900.009E+07
+ alfav           = 000.000E+07
+ alqav           = 100.001E+07
+ alkav           = 200.002E+07
+ rbi0            = 300.003E+07
+ rbx             = 400.004E+07
+ fgeo            = 500.005E+07
+ fdqr0           = 600.006E+07
+ fcrbi           = 700.007E+07
+ fqi             = 800.008E+07
+ re              = 900.009E+07
+ rcx             = 000.000E+07
+ itss            = 100.001E+07
+ msf             = 200.002E+07
+ iscs            = 300.003E+07
+ msc             = 400.004E+07
+ tsf             = 500.005E+07
+ rsu             = 600.006E+07
+ csu             = 700.007E+07
+ cjei0           = 800.008E+07
+ vdei            = 900.009E+07
+ zei             = 000.000E+07
+ ajei            = 100.001E+07
*aljei
+ cjep0           = 200.002E+07
+ vdep            = 300.003E+07
+ zep             = 400.004E+07
+ ajep            = 500.005E+07
*aljep
+ cjci0           = 600.006E+07
+ vdci            = 700.007E+07
+ zci             = 800.008E+07
+ vptci           = 900.009E+07
+ cjcx0           = 000.000E+07
+ vdcx            = 100.001E+07
+ zcx             = 200.002E+07
+ vptcx           = 300.003E+07
+ fbcpar          = 400.004E+07
*+ fbc
+ fbepar          = 500.005E+07
*+ fbe
+ cjs0            = 600.006E+07
+ vds             = 700.007E+07
+ zs              = 800.008E+07
+ vpts            = 900.009E+07
+ cscp0           = 000.000E+07
+ vdsp            = 100.001E+07
+ zsp             = 200.002E+07
+ vptsp           = 300.003E+07
+ t0              = 400.004E+07
+ dt0h            = 500.005E+07
+ tbvl            = 600.006E+07
+ tef0            = 700.007E+07
+ gtfe            = 800.008E+07
+ thcs            = 900.009E+07
+ ahc             = 000.000E+07
*alhc
+ fthc            = 100.001E+07
+ rci0            = 200.002E+07
+ vlim            = 300.003E+07
+ vces            = 400.004E+07
+ vpt             = 500.005E+07
+ aick            = 600.006E+07
+ delck           = 700.007E+07
+ tr              = 800.008E+07
+ vcbar           = 900.009E+07
+ icbar           = 000.000E+07
+ acbar           = 100.001E+07
+ cbepar          = 200.002E+07
*ceox
+ cbcpar          = 300.003E+07
*ccox
+ alqf            = 400.004E+07
+ alit            = 500.005E+07
+ flnqs           = 6
+ kf              = 700.007E+07
+ af              = 800.008E+07
+ cfbe            = 9
+ flcono          = 0
+ kfre            = 100.001E+07
+ afre            = 200.002E+07
+ latb            = 300.003E+07
+ latl            = 400.004E+07
+ vgb             = 500.005E+07
+ alt0            = 600.006E+07
+ kt0             = 700.007E+07
+ zetaci          = 800.008E+07
+ alvs            = 900.009E+07
+ alces           = 000.000E+07
+ zetarbi         = 100.001E+07
+ zetarbx         = 200.002E+07
+ zetarcx         = 300.003E+07
+ zetare          = 400.004E+07
+ zetacx          = 500.005E+07
+ vge             = 600.006E+07
+ vgc             = 700.007E+07
+ vgs             = 800.008E+07
+ f1vg            = 900.009E+07
+ f2vg            = 000.000E+07
+ zetact          = 100.001E+07
+ zetabet         = 200.002E+07
+ alb             = 300.003E+07
+ dvgbe           = 400.004E+07
+ zetahjei        = 500.005E+07
+ zetavgbe        = 600.006E+07
+ flsh            = 7
+ rth             = 800.008E+07
+ zetarth         = 900.009E+07
+ alrth           = 000.000E+07
+ cth             = 100.001E+07
+ flcomp          = 200.002E+07
+ vbe_max         = 300.003E+07
+ vbc_max         = 400.004E+07
+ vce_max         = 500.005E+07
+)

* LTspice Gummel-Poon parameters.
.MODEL _6_NPN_GUMMELPOON NPN(  
+     IS=000.000E+07
+     NF=100.001E+07
+     ISE=200.002E+07
+     NE=300.003E+07
+     BF=400.004E+07
+     IKF=500.005E+07
+     VAF=600.006E+07
+     NR=700.007E+07
+     ISC=800.008E+07
+     NC=900.009E+07
*
+     BVCBO=1
+     NBVCBO=2
+     TBVCBO1=3
+     TBVCBO2=4
+     BVBE=5
+     IBVBE=6
+     NBVBE=7
+)

* AKO model.
.MODEL _7_NPN_GUMMELPOON AKO:_6_NPN_GUMMELPOON
