* EESchema Netlist Version 1.0 (Spice format) creation date: 26/11/2005-21:12:08

.AC 10 1Meg *1.2

R12  1 3 22K
R11  2 3 100
L1  3 1 100mH
R10  5 4 220
C3  5 0 10uF
C2  9 0 1nF
R8  4 0 2.2K
Q3  1 9 4 4 Q2N2222
V2  8 0 AC 0.1
C1  11 8 1UF
V1  2 0 DC 12V
R2  11 0 10K
R6  2 11 22K
R5  2 12 22K
R1  12 0 10K
R7  7 0 470
R4  2 9 1K
R3  2 10 1K
Q2  9 12 7 7 Q2N2222
Q1  10 11 7 7 Q2N2222

.plot ac v(nodes) (-1,5)

.end
