.title KiCad schematic
.include "opamp.lib"
.save all
.probe alli
.tran 10u 10m

V3 GND Net-_U1-V-_ ( 5 ) 
R2 Net-_U1--_ Net-_R2-Pad2_ 10k 
XU1 Net-_U1-+_ Net-_U1--_ Net-_U1-V+_ Net-_U1-V-_ Net-_R2-Pad2_ uopamp_lvl2 
V2 Net-_U1-V+_ GND ( 5 ) 
V1 Net-_U1-+_ GND SIN( 0 100m 1k    ) 
R1 GND Net-_U1--_ 10k 
.end
