*
* bjts.lib.spice
* 

* All parameter values are made up and physically nonsensical.
* Commented out some parameters to avoid making test code overly long.

* First, Gummel-Poon.

*
.MODEL _0_NPN_GUMMELPOON NPN(  
+     IS=000.000E+07
+     NF=100.001E+07
+     ISE=200.002E+07
+     NE=300.003E+07
+     BF=400.004E+07
+     IKF=500.005E+07
+     VAF=600.006E+07
+     NR=700.007E+07
+     ISC=800.008E+07
+     NC=900.009E+07
+)
*+     BR=1.111E-05 
*+     IKR=2.222E-04 
*+     VAR=3.333E-03 
*+     RB=4.444E-02  
*+     IRB=5.555E-01 
*+     RBM=6.666E-00    
*+     RE=7.777E*+01 
*+     RC=8.888E*+02
*+     XTB=9.999E*+03  
*+     EG=0.000E*+04 
*+     XTI=1.111E*+05 
*+     CJE=2.222E*+06 
*+     VJE=3.333E*+07 
*+     MJE=4.444E*+08 
*+     TF=5.555E*+09 
*+     XTF=6.666E*+10 
*+     VTF=7.777E*+11   
*+     ITF=8.888E*+12 
*+     PTF=9.999E*+13  
*+     CJC=0.000E*+14 
*+     VJC=1.111E*+15 
*+     MJC=2.2222   
*+     XCJC=3.3333 
*+     TR=4.4444
*+     CJS=5.5555 
*+     VJS=6.6666 
*+     MJS=7.7777
*+     FC=8.8888 ) 
* 

*
.MODEL _1_PNP_GUMMELPOON PNP( level = 1. ; Decimal separator must be accepted too.
+     IS=000.000E+07
+     NF=100.001E+07
+     ISE=200.002E+07
+     NE=300.003E+07
+     BF=400.004E+07
+     IKF=500.005E+07
+     VAF=600.006E+07
+     NR=700.007E+07
+     ISC=800.008E+07
+     NC=900.009E+07
+)
*+     BR=1.111E-05 
*+     IKR=2.222E-04 
*+     VAR=3.333E-03 
*+     RB=4.444E-02  
*+     IRB=5.555E-01 
*+     RBM=6.666E-00    
*+     RE=7.777E*+01 
*+     RC=8.888E*+02
*+     XTB=9.999E*+03  
*+     EG=0.000E*+04 
*+     XTI=1.111E*+05 
*+     CJE=2.222E*+06 
*+     VJE=3.333E*+07 
*+     MJE=4.444E*+08 
*+     TF=5.555E*+09 
*+     XTF=6.666E*+10 
*+     VTF=7.777E*+11   
*+     ITF=8.888E*+12 
*+     PTF=9.999E*+13  
*+     CJC=0.000E*+14 
*+     VJC=1.111E*+15 
*+     MJC=2.2222   
*+     XCJC=3.3333 
*+     TR=4.4444
*+     CJS=5.5555 
*+     VJS=6.6666 
*+     MJS=7.7777
*+     FC=8.8888 ) 
* 


* VBIC.

.model _2_NPN_VBIC NPN( level=4
+ rcx             = 000.000E+07
+ rci             = 100.001E+07
+ vo              = 200.002E+07
+ gamm            = 300.003E+07
+ hrcf            = 400.004E+07
+ rbx             = 500.005E+07
+ rbi             = 600.006E+07
+ re              = 700.007E+07
+ rs              = 800.008E+07
+ rbp             = 900.009E+07
+)
*+ is              = 123.456E+07
*+ nf              = 123.456E+07
*+ nr              = 123.456E+07
*+ fc              = 123.456E+07
*+ cbeo            = 123.456E+07
*+ cje             = 123.456E+07
*+ pe              = 123.456E+07
*+ me              = 123.456E+07
*+ aje             = 123.456E+07
*+ cbco            = 123.456E+07
*+ cjc             = 123.456E+07
*+ qco             = 123.456E+07
*+ cjep            = 123.456E+07
*+ pc              = 123.456E+07
*+ mc              = 123.456E+07
*+ ajc             = 123.456E+07
*+ cjcp            = 123.456E+07
*+ ps              = 123.456E+07
*+ ms              = 123.456E+07
*+ ajs             = 123.456E+07
*+ ibei            = 123.456E+07
*+ wbe             = 123.456E+07
*+ nei             = 123.456E+07
*+ iben            = 123.456E+07
*+ nen             = 123.456E+07
*+ ibci            = 123.456E+07
*+ nci             = 123.456E+07
*+ ibcn            = 123.456E+07
*+ ncn             = 123.456E+07
*+ avc1            = 123.456E+07
*+ avc2            = 123.456E+07
*+ isp             = 123.456E+07
*+ wsp             = 123.456E+07
*+ nfp             = 123.456E+07
*+ ibeip           = 123.456E+07
*+ ibenp           = 123.456E+07
*+ ibcip           = 123.456E+07
*+ ncip            = 123.456E+07
*+ ibcnp           = 123.456E+07
*+ ncnp            = 123.456E+07
*+ vef             = 123.456E+07
*+ ver             = 123.456E+07
*+ ikf             = 123.456E+07
*+ ikr             = 123.456E+07
*+ ikp             = 123.456E+07
*+ tf              = 123.456E+07
*+ qtf             = 123.456E+07
*+ xtf             = 123.456E+07
*+ vtf             = 123.456E+07
*+ itf             = 123.456E+07
*+ tr              = 123.456E+07
*+ td              = 123.456E+07
*+ kfn             = 123.456E+07
*+ afn             = 123.456E+07
*+ bfn             = 123.456E+07
*+ xre             = 123.456E+07
*+ xrb             = 123.456E+07
*+ xrbi            = 123.456E+07
*+ xrc             = 123.456E+07
*+ xrci            = 123.456E+07
*+ xrs             = 123.456E+07
*+ xvo             = 123.456E+07
*+ ea              = 123.456E+07
*+ eaie            = 123.456E+07
*+ eaic            = 123.456E+07
*+ eais            = 123.456E+07
*+ eane            = 123.456E+07
*+ eanc            = 123.456E+07
*+ eans            = 123.456E+07
*+ xis             = 123.456E+07
*+ xii             = 123.456E+07
*+ xin             = 123.456E+07
*+ tnf             = 123.456E+07
*+ tavc            = 123.456E+07
*+ rth             = 123.456E+07
*+ cth             = 123.456E+07
*+ vrt             = 123.456E+07
*+ art             = 123.456E+07
*+ ccso            = 123.456E+07
*+ qbm             = 123.456E+07
*+ nkf             = 123.456E+07
*+ xikf            = 123.456E+07
*+ xrcx            = 123.456E+07
*+ xrbx            = 123.456E+07
*+ xrbp            = 123.456E+07
*+ isrr            = 123.456E+07
*+ xisr            = 123.456E+07
*+ dear            = 123.456E+07
*+ eap             = 123.456E+07
*+ vbbe            = 123.456E+07
*+ nbbe            = 123.456E+07
*+ ibbe            = 123.456E+07
*+ tvbbe1          = 123.456E+07
*+ tvbbe2          = 123.456E+07
*+ tnbbe           = 123.456E+07
*+ ebbe            = 123.456E+07
*+ dtemp           = 123.456E+07
*+ vers            = 123.456E+07
*+ vref            = 123.456E+07
*+ vbe_max         = 123.456E+07
*+ vbc_max         = 123.456E+07
*+ vce_max         = 123.456E+07
*+)

.model _3_PNP_VBIC PNP( level=4.0
+ rcx             = 000.000E+07
+ rci             = 100.001E+07
+ vo              = 200.002E+07
+ gamm            = 300.003E+07
+ hrcf            = 400.004E+07
+ rbx             = 500.005E+07
+ rbi             = 600.006E+07
+ re              = 700.007E+07
+ rs              = 800.008E+07
+ rbp             = 900.009E+07
+)
*+ is              = 123.456E+07
*+ nf              = 123.456E+07
*+ nr              = 123.456E+07
*+ fc              = 123.456E+07
*+ cbeo            = 123.456E+07
*+ cje             = 123.456E+07
*+ pe              = 123.456E+07
*+ me              = 123.456E+07
*+ aje             = 123.456E+07
*+ cbco            = 123.456E+07
*+ cjc             = 123.456E+07
*+ qco             = 123.456E+07
*+ cjep            = 123.456E+07
*+ pc              = 123.456E+07
*+ mc              = 123.456E+07
*+ ajc             = 123.456E+07
*+ cjcp            = 123.456E+07
*+ ps              = 123.456E+07
*+ ms              = 123.456E+07
*+ ajs             = 123.456E+07
*+ ibei            = 123.456E+07
*+ wbe             = 123.456E+07
*+ nei             = 123.456E+07
*+ iben            = 123.456E+07
*+ nen             = 123.456E+07
*+ ibci            = 123.456E+07
*+ nci             = 123.456E+07
*+ ibcn            = 123.456E+07
*+ ncn             = 123.456E+07
*+ avc1            = 123.456E+07
*+ avc2            = 123.456E+07
*+ isp             = 123.456E+07
*+ wsp             = 123.456E+07
*+ nfp             = 123.456E+07
*+ ibeip           = 123.456E+07
*+ ibenp           = 123.456E+07
*+ ibcip           = 123.456E+07
*+ ncip            = 123.456E+07
*+ ibcnp           = 123.456E+07
*+ ncnp            = 123.456E+07
*+ vef             = 123.456E+07
*+ ver             = 123.456E+07
*+ ikf             = 123.456E+07
*+ ikr             = 123.456E+07
*+ ikp             = 123.456E+07
*+ tf              = 123.456E+07
*+ qtf             = 123.456E+07
*+ xtf             = 123.456E+07
*+ vtf             = 123.456E+07
*+ itf             = 123.456E+07
*+ tr              = 123.456E+07
*+ td              = 123.456E+07
*+ kfn             = 123.456E+07
*+ afn             = 123.456E+07
*+ bfn             = 123.456E+07
*+ xre             = 123.456E+07
*+ xrb             = 123.456E+07
*+ xrbi            = 123.456E+07
*+ xrc             = 123.456E+07
*+ xrci            = 123.456E+07
*+ xrs             = 123.456E+07
*+ xvo             = 123.456E+07
*+ ea              = 123.456E+07
*+ eaie            = 123.456E+07
*+ eaic            = 123.456E+07
*+ eais            = 123.456E+07
*+ eane            = 123.456E+07
*+ eanc            = 123.456E+07
*+ eans            = 123.456E+07
*+ xis             = 123.456E+07
*+ xii             = 123.456E+07
*+ xin             = 123.456E+07
*+ tnf             = 123.456E+07
*+ tavc            = 123.456E+07
*+ rth             = 123.456E+07
*+ cth             = 123.456E+07
*+ vrt             = 123.456E+07
*+ art             = 123.456E+07
*+ ccso            = 123.456E+07
*+ qbm             = 123.456E+07
*+ nkf             = 123.456E+07
*+ xikf            = 123.456E+07
*+ xrcx            = 123.456E+07
*+ xrbx            = 123.456E+07
*+ xrbp            = 123.456E+07
*+ isrr            = 123.456E+07
*+ xisr            = 123.456E+07
*+ dear            = 123.456E+07
*+ eap             = 123.456E+07
*+ vbbe            = 123.456E+07
*+ nbbe            = 123.456E+07
*+ ibbe            = 123.456E+07
*+ tvbbe1          = 123.456E+07
*+ tvbbe2          = 123.456E+07
*+ tnbbe           = 123.456E+07
*+ ebbe            = 123.456E+07
*+ dtemp           = 123.456E+07
*+ vers            = 123.456E+07
*+ vref            = 123.456E+07
*+ vbe_max         = 123.456E+07
*+ vbc_max         = 123.456E+07
*+ vce_max         = 123.456E+07
*+)


* HICUM/L2

.model _4_NPN_HICUML2 NPN( level=8.00
+ c10             = 000.000E+07
+ qp0             = 100.001E+07
+ ich             = 200.002E+07
+ hf0             = 300.003E+07
+ hfe             = 400.004E+07
+ hfc             = 500.005E+07
+ hjei            = 600.006E+07
+ ahjei           = 700.007E+07
+ rhjei           = 800.008E+07
+ hjci            = 900.009E+07
+)
*+ ibeis           = 123.456E+07
*+ mbei            = 123.456E+07
*+ ireis           = 123.456E+07
*+ mrei            = 123.456E+07
*+ ibeps           = 123.456E+07
*+ mbep            = 123.456E+07
*+ ireps           = 123.456E+07
*+ mrep            = 123.456E+07
*+ mcf             = 123.456E+07
*+ tbhrec          = 123.456E+07
*+ ibcis           = 123.456E+07
*+ mbci            = 123.456E+07
*+ ibcxs           = 123.456E+07
*+ mbcx            = 123.456E+07
*+ ibets           = 123.456E+07
*+ abet            = 123.456E+07
*+ tunode          = 123.456E+07
*+ favl            = 123.456E+07
*+ qavl            = 123.456E+07
*+ kavl            = 123.456E+07
*+ alfav           = 123.456E+07
*+ alqav           = 123.456E+07
*+ alkav           = 123.456E+07
*+ rbi0            = 123.456E+07
*+ rbx             = 123.456E+07
*+ fgeo            = 123.456E+07
*+ fdqr0           = 123.456E+07
*+ fcrbi           = 123.456E+07
*+ fqi             = 123.456E+07
*+ re              = 123.456E+07
*+ rcx             = 123.456E+07
*+ itss            = 123.456E+07
*+ msf             = 123.456E+07
*+ iscs            = 123.456E+07
*+ msc             = 123.456E+07
*+ tsf             = 123.456E+07
*+ rsu             = 123.456E+07
*+ csu             = 123.456E+07
*+ cjei0           = 123.456E+07
*+ vdei            = 123.456E+07
*+ zei             = 123.456E+07
*+ ajei            = 123.456E+07
*+ aljei           = 123.456E+07
*+ cjep0           = 123.456E+07
*+ vdep            = 123.456E+07
*+ zep             = 123.456E+07
*+ ajep            = 123.456E+07
*+ aljep           = 123.456E+07
*+ cjci0           = 123.456E+07
*+ vdci            = 123.456E+07
*+ zci             = 123.456E+07
*+ vptci           = 123.456E+07
*+ cjcx0           = 123.456E+07
*+ vdcx            = 123.456E+07
*+ zcx             = 123.456E+07
*+ vptcx           = 123.456E+07
*+ fbcpar          = 123.456E+07
*+ fbc             = 123.456E+07
*+ fbepar          = 123.456E+07
*+ fbe             = 123.456E+07
*+ cjs0            = 123.456E+07
*+ vds             = 123.456E+07
*+ zs              = 123.456E+07
*+ vpts            = 123.456E+07
*+ cscp0           = 123.456E+07
*+ vdsp            = 123.456E+07
*+ zsp             = 123.456E+07
*+ vptsp           = 123.456E+07
*+ t0              = 123.456E+07
*+ dt0h            = 123.456E+07
*+ tbvl            = 123.456E+07
*+ tef0            = 123.456E+07
*+ gtfe            = 123.456E+07
*+ thcs            = 123.456E+07
*+ ahc             = 123.456E+07
*+ alhc            = 123.456E+07
*+ fthc            = 123.456E+07
*+ rci0            = 123.456E+07
*+ vlim            = 123.456E+07
*+ vces            = 123.456E+07
*+ vpt             = 123.456E+07
*+ aick            = 123.456E+07
*+ delck           = 123.456E+07
*+ tr              = 123.456E+07
*+ vcbar           = 123.456E+07
*+ icbar           = 123.456E+07
*+ acbar           = 123.456E+07
*+ cbepar          = 123.456E+07
*+ ceox            = 123.456E+07
*+ cbcpar          = 123.456E+07
*+ ccox            = 123.456E+07
*+ alqf            = 123.456E+07
*+ alit            = 123.456E+07
*+ flnqs           = 123.456E+07
*+ kf              = 123.456E+07
*+ af              = 123.456E+07
*+ cfbe            = 123.456E+07
*+ flcono          = 123.456E+07
*+ kfre            = 123.456E+07
*+ afre            = 123.456E+07
*+ latb            = 123.456E+07
*+ latl            = 123.456E+07
*+ vgb             = 123.456E+07
*+ alt0            = 123.456E+07
*+ kt0             = 123.456E+07
*+ zetaci          = 123.456E+07
*+ alvs            = 123.456E+07
*+ alces           = 123.456E+07
*+ zetarbi         = 123.456E+07
*+ zetarbx         = 123.456E+07
*+ zetarcx         = 123.456E+07
*+ zetare          = 123.456E+07
*+ zetacx          = 123.456E+07
*+ vge             = 123.456E+07
*+ vgc             = 123.456E+07
*+ vgs             = 123.456E+07
*+ f1vg            = 123.456E+07
*+ f2vg            = 123.456E+07
*+ zetact          = 123.456E+07
*+ zetabet         = 123.456E+07
*+ alb             = 123.456E+07
*+ dvgbe           = 123.456E+07
*+ zetahjei        = 123.456E+07
*+ zetavgbe        = 123.456E+07
*+ flsh            = 123.456E+07
*+ rth             = 123.456E+07
*+ zetarth         = 123.456E+07
*+ alrth           = 123.456E+07
*+ cth             = 123.456E+07
*+ flcomp          = 123.456E+07
*+ vbe_max         = 123.456E+07
*+ vbc_max         = 123.456E+07
*+ vce_max         = 123.456E+07
*+)

.model _5_PNP_HICUML2 PNP( level=8
+ c10             = 000.000E+07
+ qp0             = 100.001E+07
+ ich             = 200.002E+07
+ hf0             = 300.003E+07
+ hfe             = 400.004E+07
+ hfc             = 500.005E+07
+ hjei            = 600.006E+07
+ ahjei           = 700.007E+07
+ rhjei           = 800.008E+07
+ hjci            = 900.009E+07
+)
*+ ibeis           = 123.456E+07
*+ mbei            = 123.456E+07
*+ ireis           = 123.456E+07
*+ mrei            = 123.456E+07
*+ ibeps           = 123.456E+07
*+ mbep            = 123.456E+07
*+ ireps           = 123.456E+07
*+ mrep            = 123.456E+07
*+ mcf             = 123.456E+07
*+ tbhrec          = 123.456E+07
*+ ibcis           = 123.456E+07
*+ mbci            = 123.456E+07
*+ ibcxs           = 123.456E+07
*+ mbcx            = 123.456E+07
*+ ibets           = 123.456E+07
*+ abet            = 123.456E+07
*+ tunode          = 123.456E+07
*+ favl            = 123.456E+07
*+ qavl            = 123.456E+07
*+ kavl            = 123.456E+07
*+ alfav           = 123.456E+07
*+ alqav           = 123.456E+07
*+ alkav           = 123.456E+07
*+ rbi0            = 123.456E+07
*+ rbx             = 123.456E+07
*+ fgeo            = 123.456E+07
*+ fdqr0           = 123.456E+07
*+ fcrbi           = 123.456E+07
*+ fqi             = 123.456E+07
*+ re              = 123.456E+07
*+ rcx             = 123.456E+07
*+ itss            = 123.456E+07
*+ msf             = 123.456E+07
*+ iscs            = 123.456E+07
*+ msc             = 123.456E+07
*+ tsf             = 123.456E+07
*+ rsu             = 123.456E+07
*+ csu             = 123.456E+07
*+ cjei0           = 123.456E+07
*+ vdei            = 123.456E+07
*+ zei             = 123.456E+07
*+ ajei            = 123.456E+07
*+ aljei           = 123.456E+07
*+ cjep0           = 123.456E+07
*+ vdep            = 123.456E+07
*+ zep             = 123.456E+07
*+ ajep            = 123.456E+07
*+ aljep           = 123.456E+07
*+ cjci0           = 123.456E+07
*+ vdci            = 123.456E+07
*+ zci             = 123.456E+07
*+ vptci           = 123.456E+07
*+ cjcx0           = 123.456E+07
*+ vdcx            = 123.456E+07
*+ zcx             = 123.456E+07
*+ vptcx           = 123.456E+07
*+ fbcpar          = 123.456E+07
*+ fbc             = 123.456E+07
*+ fbepar          = 123.456E+07
*+ fbe             = 123.456E+07
*+ cjs0            = 123.456E+07
*+ vds             = 123.456E+07
*+ zs              = 123.456E+07
*+ vpts            = 123.456E+07
*+ cscp0           = 123.456E+07
*+ vdsp            = 123.456E+07
*+ zsp             = 123.456E+07
*+ vptsp           = 123.456E+07
*+ t0              = 123.456E+07
*+ dt0h            = 123.456E+07
*+ tbvl            = 123.456E+07
*+ tef0            = 123.456E+07
*+ gtfe            = 123.456E+07
*+ thcs            = 123.456E+07
*+ ahc             = 123.456E+07
*+ alhc            = 123.456E+07
*+ fthc            = 123.456E+07
*+ rci0            = 123.456E+07
*+ vlim            = 123.456E+07
*+ vces            = 123.456E+07
*+ vpt             = 123.456E+07
*+ aick            = 123.456E+07
*+ delck           = 123.456E+07
*+ tr              = 123.456E+07
*+ vcbar           = 123.456E+07
*+ icbar           = 123.456E+07
*+ acbar           = 123.456E+07
*+ cbepar          = 123.456E+07
*+ ceox            = 123.456E+07
*+ cbcpar          = 123.456E+07
*+ ccox            = 123.456E+07
*+ alqf            = 123.456E+07
*+ alit            = 123.456E+07
*+ flnqs           = 123.456E+07
*+ kf              = 123.456E+07
*+ af              = 123.456E+07
*+ cfbe            = 123.456E+07
*+ flcono          = 123.456E+07
*+ kfre            = 123.456E+07
*+ afre            = 123.456E+07
*+ latb            = 123.456E+07
*+ latl            = 123.456E+07
*+ vgb             = 123.456E+07
*+ alt0            = 123.456E+07
*+ kt0             = 123.456E+07
*+ zetaci          = 123.456E+07
*+ alvs            = 123.456E+07
*+ alces           = 123.456E+07
*+ zetarbi         = 123.456E+07
*+ zetarbx         = 123.456E+07
*+ zetarcx         = 123.456E+07
*+ zetare          = 123.456E+07
*+ zetacx          = 123.456E+07
*+ vge             = 123.456E+07
*+ vgc             = 123.456E+07
*+ vgs             = 123.456E+07
*+ f1vg            = 123.456E+07
*+ f2vg            = 123.456E+07
*+ zetact          = 123.456E+07
*+ zetabet         = 123.456E+07
*+ alb             = 123.456E+07
*+ dvgbe           = 123.456E+07
*+ zetahjei        = 123.456E+07
*+ zetavgbe        = 123.456E+07
*+ flsh            = 123.456E+07
*+ rth             = 123.456E+07
*+ zetarth         = 123.456E+07
*+ alrth           = 123.456E+07
*+ cth             = 123.456E+07
*+ flcomp          = 123.456E+07
*+ vbe_max         = 123.456E+07
*+ vbc_max         = 123.456E+07
*+ vce_max         = 123.456E+07
*+)
