* EESchema Netlist Version 1.1 (Spice format) creation date: 05/01/2014 19:00:38

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
R12  /VOUT Net-_L1-Pad1_ 22K		
R11  +12V Net-_L1-Pad1_ 100		
L1  Net-_L1-Pad1_ /VOUT 100mH		
R10  Net-_C3-Pad1_ Net-_Q3-Pad3_ 220		
C3  Net-_C3-Pad1_ 0 10uF		
C2  Net-_C2-Pad1_ 0 1nF		
R8  Net-_Q3-Pad3_ 0 2.2K		
Q3  /VOUT Net-_C2-Pad1_ Net-_Q3-Pad3_ Net-_Q3-Pad3_ Q2N2222		
V2  Net-_C1-Pad2_ 0 AC 0.1		
C1  /VIN Net-_C1-Pad2_ 1UF		
V1  +12V 0 DC 12V		
R2  /VIN 0 10K		
R6  +12V /VIN 22K		
R5  +12V Net-_Q2-Pad2_ 22K		
R1  Net-_Q2-Pad2_ 0 10K		
R7  Net-_Q1-Pad3_ 0 470		
R4  +12V Net-_C2-Pad1_ 1K		
R3  +12V Net-_Q1-Pad1_ 1K		
Q2  Net-_C2-Pad1_ Net-_Q2-Pad2_ Net-_Q1-Pad3_ Net-_Q1-Pad3_ Q2N2222		
Q1  Net-_Q1-Pad1_ /VIN Net-_Q1-Pad3_ Net-_Q1-Pad3_ Q2N2222		

.model Q2N2222 npn (bf=200)
.print tran v(nodes)
.print dc v(nodes)
.tran 10 10000 10 > pspice.dat

.end
